----------------------------------------------------------------------------------
-- Autor: 			Marcel Cholodecki
-- Numer albumu: 	275818
-- Projekt:			Gra kolko i krzyzyk
--
-- Pakiet:			my_package.vhd
-- Opis:				Typy wykorzystane w projekcie
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package my_package is

	-- Typ wyliczeniowy do obslugi stanu planszy
	type GAME_t is ('-', 'O', 'X');
	type GAME_t_Vector is ARRAY (8 downto 0) of GAME_t;

end my_package;

package body my_package is
end my_package;
