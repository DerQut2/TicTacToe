----------------------------------------------------------------------------------
-- Autor: 			Marcel Cholodecki
-- Numer albumu: 	275818
-- Projekt:			Gra kolko i krzyzyk
--
-- Pakiet:			my_package.vhd
-- Opis:				Typy wyliczeniowe wykorzystane w projekcie
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package my_package is

	-- Typ wyliczeniowy do obslugi stanu planszy
	type gametype is ('X', 'O', '-');

end my_package;

package body my_package is
end my_package;
